event Ev1 is {informal #ErrorOverflowMailBox# }
event Ev is {send sample to {moteur}0}
event Ev3 is { send sample to {moteur}0}
event Ev4 is { receive sample from any}
event Ev5 is {receive sample from any}
event Debut is {send debut to {moteur}0}
event Sample is {send sample to {moteur}0}
event Sample2 is { send sample to {moteur}0}
event sample3 is {send sample to {moteur}0}
event send2 is { send avance to {moteur}0}
event ack1 is { receive OK from any}
event ack2 is { receive OK from any}

event Fin is { send fin to {moteur}0}

cdl Exemple9 is {
	main is { SEQniveau1 || SEQniveau2 || SEQniveau3 }
}

activity SEQniveau1 is {
	event Debut; event Sample2; event sample3;
	{ 
		loop 3 event Sample2
	[]	{
			event sample3; 
			{
				event ack1  
			[]	event ack2
			}
		}
	}
}

activity SEQniveau2 is {
	event Ev;
	{ 
		loop 3 event Ev
	[]	event ack1 
	[]	
		{
			event Ev3  
		[]	event Ev4
		[]	{ event Sample; event Ev5 } 
		}
	}
}

activity SEQniveau3 is {
	event Debut; event Fin
}


