activity HMI0_login is {
	event {send t_msg {id = 0, body = t_body.login(true)} to {SM}1}
}

activity HMI1_login is {
	event {send t_msg {id = 1, body = t_body.login(true)} to {SM}1}
}

activity HMI2_login is {
	event {send t_msg {id = 2, body = t_body.login(true)} to {SM}1}
[]	event {send t_msg {id = 2, body = t_body.login(false)} to {SM}1}
}

activity HMI0_logout is {
	event {send t_msg {id = 0, body = t_body.logout} to {SM}1}
}

activity HMI1_logout is {
	event {send t_msg {id = 1, body = t_body.logout} to {SM}1}
}

activity HMI2_logout is {
	event {send t_msg {id = 2, body = t_body.logout} to {SM}1}
}

activity HMI0_operate is {
	event {send t_msg {id = 0, body = t_body.operate} to {SM}1}
}

activity HMI1_operate is {
	event {send t_msg {id = 1, body = t_body.operate} to {SM}1}
}

activity HMI2_operate is {
	event {send t_msg {id = 2, body = t_body.operate} to {SM}1}
}

activity HMI0_login_and_logout is {
	HMI0_login;
	HMI0_logout
}

activity HMI1_login_and_logout is {
	HMI1_login;
	HMI1_logout
}

activity HMI2_login_and_logout is {
	HMI2_login;
	HMI2_logout
}

activity HMI0_login_operate_and_logout is {
	HMI0_login;
	HMI0_operate;
	HMI0_logout
}

activity HMI1_login_operate_and_logout is {
	HMI1_login;
	HMI1_operate;
	HMI1_logout
}

activity HMI2_login_operate_and_logout is {
	HMI2_login;
	HMI2_operate;
	HMI2_logout
}

event ack_HMI0 is {receive t_msg {id = 0, body = t_body.ack(true)} from {SM}1}
event nack_HMI0 is {receive t_msg {id = 0, body = t_body.ack(false)} from {SM}1}
event ack_HMI1 is {receive t_msg {id = 1, body = t_body.ack(true)} from {SM}1}
event nack_HMI1 is {receive t_msg {id = 1, body = t_body.ack(false)} from {SM}1}
event ack_HMI2 is {receive t_msg {id = 2, body = t_body.ack(true)} from {SM}1}
event nack_HMI2 is {receive t_msg {id = 2, body = t_body.ack(false)} from {SM}1}

property HMI0_is_right is {
	start -- / / nack_HMI0 / -> reject
}

property HMI1_is_right is {
	start -- / / nack_HMI1 / -> reject
}

property HMI2_is_wrong is {
	start -- / / nack_HMI2 / -> success
}

event any_login is {receive t_msg {id = any, body = t_body.login(any)} from {env}1 to {SM}1}
event any_ack is {send t_msg {id = any, body = t_body.ack(any)} from {SM}1 to {env}1}

property matches_any_login is {
	start -- / / any_login / -> success
}

property matches_any_ack is {
	start -- / / any_ack / -> success
}

property ack_follows_login is {
	start -- / / any_login / -> wait;
	wait -- / / any_ack / -> start;
	wait -- / / / -> reject
}

cdl empty is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		skip
	}
}

cdl HMI0_login is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login
	}
}

cdl HMI0_login_and_logout is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login_and_logout
	}
}

cdl HMI0_login_operate_and_logout is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login_operate_and_logout
	}
}

cdl HMI0n1_login is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login
	||	HMI1_login
	}
}

cdl HMI0n1_login_and_logout is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login_and_logout
	||  HMI1_login_and_logout
	}
}

cdl HMI0n1_login_operate_and_logout is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login_operate_and_logout
	||	HMI1_login_operate_and_logout
	}
}

cdl HMI0n2_login is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login
	||	HMI2_login
	}
}

cdl HMI0n2_login_and_logout is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login_and_logout
	||  HMI2_login_and_logout
	}
}

cdl HMI0n2_login_operate_and_logout is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login_operate_and_logout
	||	HMI2_login_operate_and_logout
	}
}

cdl HMI0n1n2_login is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login
	||	HMI1_login
	||	HMI2_login
	}
}

cdl HMI0n1n2_login_and_logout is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login_and_logout
	||  HMI1_login_and_logout
	||  HMI2_login_and_logout
	}
}

cdl HMI0n1n2_login_operate_and_logout is {
	properties
		HMI0_is_right,
		HMI1_is_right,
		HMI2_is_wrong,
		matches_any_login,
		matches_any_ack,
		ack_follows_login

	main is {
		HMI0_login_operate_and_logout
	||	HMI1_login_operate_and_logout
	||	HMI2_login_operate_and_logout
	}
}